package dmaRegConfigPkg;

parameter ADDRESSWIDTH = 16;
parameter DATAWIDTH = 8;
parameter CHANNELS = 4;
parameter REGISTERADDRESS = 4;

endpackage
